* Randles Circuit Model for Li-ion Battery (5-stage Cauer Warburg, ngspice-ready)
* ------------------------------------------------------------
* Top-level parameters (replace defaults or override when invoking ngspice)
.param Ru_val = 0.02     ; Ohmic Resistance (Ohm) - default
.param Rct_val = 0.05   ; Charge Transfer Resistance (Ohm)
.param Cdl_val = 0.0005   ; Double Layer Capacitance (F)
.param Wsig_val = 10 ; Warburg coefficient (Ohm) - total diffusion resistance approx
.param Tw_val = 10       ; Warburg diffusion time constant (s)



* -------------------------
* Warburg subcircuit (5-stage Cauer ladder approximating finite Warburg)
* Pins: P = input node, N = reference/ground
.subckt Warburg P N
* number of ladder stages (adjust if needed)
.param N_stages = 5

* total diffusion resistance and capacitance for the Warburg approximation
* Rw_total is taken from Wsig_val (user-supplied)
.param Rw_total = {Wsig_val}
* Cw_total computed from Tw_val / Rw_total (C = Tau / R)
.param Cw_total = {Tw_val / Rw_total}

* per-stage resistor and capacitor
.param R_each = {Rw_total / N_stages}
.param C_each = {Cw_total / N_stages}

* Ladder / Cauer network:
* Stage 1
R1 P 10 {R_each}
C1 10 N {C_each}

* Stage 2
R2 10 20 {R_each}
C2 20 N {C_each}

* Stage 3
R3 20 30 {R_each}
C3 30 N {C_each}

* Stage 4
R4 30 40 {R_each}
C4 40 N {C_each}

* Stage 5 (terminate diffusion path with capacitor to model finite/blocked diffusion)
R5 40 50 {R_each}
C5 50 N {C_each}

.ends Warburg

* -------------------------
* Main Randles cell subcircuit
* Pins: P = positive/input, N = reference/ground
.subckt RandlesCell P N
* Ru (ohmic), Cdl (double layer) in parallel with (Rct + Warburg)
R_u P 1 {Ru_val}
C_dl 1 N {Cdl_val}

R_ct 1 N {Rct_val}
* call Warburg subcircuit between node 2 and ground (N)
* X_warburg 2 N Warburg

.ends RandlesCell

* --- control ---


* --- control ---

* Test Circuit - Stimulus for EIS
V_source 100 0 AC 1V
X_cell 100 0 RandlesCell

* AC Analysis settings
.ac dec 10 0.001 10000000.0

.control
  run
  set units = si
  
  * Define the Frequency vector
  let freq = frequency
  
  * Calculate Complex Impedance
  * Note: I(V_source) is negative convention in SPICE, so we use -I to get positive Z
  let Z = V(100) / -I(V_source)
  
  * Extract Components for EIS Analysis
  let Z_mag = abs(Z)
  let Z_phase = ph(Z)
  let Z_real = real(Z)
  let Z_imag = imag(Z)
  
  * Output to console (for parsing)
  print freq Z_mag Z_phase
  
  * Save data to file
  wrdata runs/20251120034520_a0707c69/eis_data.txt Z_real Z_imag Z_mag Z_phase

.endc

.end
