
* Randles Circuit Model for Li-ion Battery

.param Ru_val = 0.02
.param Rct_val = 0.5
.param Cdl_val = 0.0005
.param Wsig_val = 0.1

.subckt Warburg P N
.param N_stages = 5

.param R_each = {Wsig_val / N_stages}
.param C_each = {N_stages / Wsig_val}

R1 P 10 {R_each}
C1 10 N {C_each}
R2 10 20 {R_each}
C2 20 N {C_each}
R3 20 30 {R_each}
C3 30 N {C_each}
R4 30 40 {R_each}
C4 40 N {C_each}
R5 40 N {R_each}
C5 40 N {C_each}
.ends

.subckt RandlesCell P N
R_u P 1 {Ru_val}       ; Ohmic resistance
C_dl 1 N {Cdl_val}     ; Double layer capacitance, in parallel with Rct+Warburg branch
R_ct 1 2 {Rct_val}     ; Charge transfer resistance
X_warburg 2 N Warburg  ; Warburg impedance in series with Rct
.ends

* exported_nodes: 1, 2, 10, 20, 30, 40, N


* --- control ---


* --- control ---

* Test Circuit - Stimulus for EIS
V_source 100 0 AC 1V
X_cell 100 0 RandlesCell

* AC Analysis settings
.ac dec 10 0.001 10000.0

.control
  run
  set units = si
  
  * Define the Frequency vector
  let freq = frequency
  
  * Calculate Complex Impedance
  * Note: I(V_source) is negative convention in SPICE, so we use -I to get positive Z
  let Z = V(100) / -I(V_source)
  
  * Extract Components for EIS Analysis
  let Z_mag = abs(Z)
  let Z_phase = ph(Z)
  let Z_real = real(Z)
  let Z_imag = imag(Z)
  
  * Output to console (for parsing)
  print freq Z_mag Z_phase
  
  * Save data to file
  wrdata runs/20251119080926_dc6af700/eis_data.txt Z_real Z_imag Z_mag Z_phase

.endc

.end
